module ram(clk, cen, wen, addr, din, dout);
	input clk;
	input cen, wen;
	input[15:0] addr; //addr[5:0] = 000000(0) ~ 111111(63)
	input[31:0] din;
	output reg[31:0] dout;
	
	reg[31:0] mem[63:0];
	
	initial
		begin
			mem[0] = 32'h0000_0000;
			mem[1] = 32'h0000_0000;
			mem[2] = 32'h0000_0000;
			mem[3] = 32'h0000_0000;
			mem[4] = 32'h0000_0000;
			mem[5] = 32'h0000_0000;
			mem[6] = 32'h0000_0000;
			mem[7] = 32'h0000_0000;
			mem[8] = 32'h0000_0000;
			mem[9] = 32'h0000_0000;
			
			mem[10] = 32'h0000_0000;
			mem[11] = 32'h0000_0000;
			mem[12] = 32'h0000_0000;
			mem[13] = 32'h0000_0000;
			mem[14] = 32'h0000_0000;
			mem[15] = 32'h0000_0000;
			mem[16] = 32'h0000_0000;
			mem[17] = 32'h0000_0000;
			mem[18] = 32'h0000_0000;
			mem[19] = 32'h0000_0000;
			
			mem[20] = 32'h0000_0000;
			mem[21] = 32'h0000_0000;
			mem[22] = 32'h0000_0000;
			mem[23] = 32'h0000_0000;
			mem[24] = 32'h0000_0000;
			mem[25] = 32'h0000_0000;
			mem[26] = 32'h0000_0000;
			mem[27] = 32'h0000_0000;
			mem[28] = 32'h0000_0000;
			mem[29] = 32'h0000_0000;
			
			mem[30] = 32'h0000_0000;
			mem[31] = 32'h0000_0000;
			mem[32] = 32'h0000_0000;
			mem[33] = 32'h0000_0000;
			mem[34] = 32'h0000_0000;
			mem[35] = 32'h0000_0000;
			mem[36] = 32'h0000_0000;
			mem[37] = 32'h0000_0000;
			mem[38] = 32'h0000_0000;
			mem[39] = 32'h0000_0000;
			
			mem[40] = 32'h0000_0000;
			mem[41] = 32'h0000_0000;
			mem[42] = 32'h0000_0000;
			mem[43] = 32'h0000_0000;
			mem[44] = 32'h0000_0000;
			mem[45] = 32'h0000_0000;
			mem[46] = 32'h0000_0000;
			mem[47] = 32'h0000_0000;
			mem[48] = 32'h0000_0000;
			mem[49] = 32'h0000_0000;
			
			mem[50] = 32'h0000_0000;
			mem[51] = 32'h0000_0000;
			mem[52] = 32'h0000_0000;
			mem[53] = 32'h0000_0000;
			mem[54] = 32'h0000_0000;
			mem[55] = 32'h0000_0000;
			mem[56] = 32'h0000_0000;
			mem[57] = 32'h0000_0000;
			mem[58] = 32'h0000_0000;
			mem[59] = 32'h0000_0000;
			
			mem[60] = 32'h0000_0000;
			mem[61] = 32'h0000_0000;
			mem[62] = 32'h0000_0000;
			mem[63] = 32'h0000_0000;
			//mem[63:0] = 0;
		end
		
	always @ (posedge clk)
		begin
			if ({cen,wen} == 2'b11)
				begin
					mem[addr[5:0]] = din; //write
					dout = 32'h0000_0000;
				end
			
			else if ({cen,wen} == 2'b10)
				begin
					dout = mem[addr[5:0]]; //read
				end
				
			else if (cen == 1'b0)
				begin
					dout = 32'h0000_0000; //meaningless output
				end
				
			else
				begin
					dout = 32'hxxxx_xxxx; //error
				end
		end
endmodule 